module char_rom (
    input  logic [6:0] ascii_addr,
    input  logic [2:0] char_row,
    output logic [7:0] data
);
    // 3-D vector to represent ascii table
    logic [7:0] char [0:127][0:7];

    initial begin
    
        // Nums
        char[7'h30] = '{
            8'b00111100,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b00111100
        };

        char[7'h31] = '{
            8'b00001000,
            8'b00011000,
            8'b00101000,
            8'b00001000,
            8'b00001000,
            8'b00001000,
            8'b00001000,
            8'b00111110
        };

        char[7'h32] = '{
            8'b00111100,
            8'b01000010,
            8'b00000010,
            8'b00000100,
            8'b00011000,
            8'b00100000,
            8'b01000000,
            8'b01111110
        };

        char[7'h33] = '{
            8'b00111100,
            8'b01000010,
            8'b00000010,
            8'b00011100,
            8'b00000010,
            8'b00000010,
            8'b01000010,
            8'b00111100
        };

        char[7'h34] = '{
            8'b00001100,
            8'b00010100,
            8'b00100100,
            8'b01000100,
            8'b01111110,
            8'b00000100,
            8'b00000100,
            8'b00000100
        };

        char[7'h35] = '{
            8'b01111110,
            8'b01000000,
            8'b01000000,
            8'b01111100,
            8'b00000010,
            8'b00000010,
            8'b01000010,
            8'b00111100
        };

        char[7'h36] = '{
            8'b00111100,
            8'b01000010,
            8'b01000000,
            8'b01111100,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b00111100
        };

        char[7'h37] = '{
            8'b01111110,
            8'b00000010,
            8'b00000100,
            8'b00000100,
            8'b00001000,
            8'b00001000,
            8'b00010000,
            8'b00010000
        };

        char[7'h38] = '{
            8'b00111100,
            8'b01000010,
            8'b01000010,
            8'b00111100,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b00111100
        };

        char[7'h39] = '{
            8'b00111100,
            8'b01000010,
            8'b01000010,
            8'b00111110,
            8'b00000010,
            8'b00000010,
            8'b01000010,
            8'b00111100
        };
        
        // Letters
        char[7'h41] = '{
            8'b00011000,
            8'b00100100,
            8'b01000010,
            8'b01000010,
            8'b01111110,
            8'b01000010,
            8'b01000010,
            8'b01000010
        };

        char[7'h42] = '{
            8'b01111100,
            8'b01000010,
            8'b01000010,
            8'b01111100,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01111100
        };

        char[7'h43] = '{
            8'b00111100,
            8'b01000010,
            8'b01000000,
            8'b01000000,
            8'b01000000,
            8'b01000000,
            8'b01000010,
            8'b00111100
        };

        char[7'h45] = '{
            8'b01111110,
            8'b01000000,
            8'b01000000,
            8'b01111100,
            8'b01000000,
            8'b01000000,
            8'b01000000,
            8'b01111110
        };

        char[7'h47] = '{
            8'b00111100,
            8'b01000010,
            8'b01000000,
            8'b01000000,
            8'b01001110,
            8'b01000010,
            8'b01000010,
            8'b00111100
        };

        char[7'h48] = '{
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01111110,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010
        };

        char[7'h49] = '{
            8'b00111100,
            8'b00011000,
            8'b00011000,
            8'b00011000,
            8'b00011000,
            8'b00011000,
            8'b00011000,
            8'b00111100
        };

        char[7'h4C] = '{
            8'b01000000,
            8'b01000000,
            8'b01000000,
            8'b01000000,
            8'b01000000,
            8'b01000000,
            8'b01000000,
            8'b01111110
        };

        char[7'h4D] = '{
            8'b01000010,
            8'b01100110,
            8'b01011010,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010
        };

        char[7'h4F] = '{
            8'b00111100,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b00111100
        };

        char[7'h50] = '{
            8'b01111100,
            8'b01000010,
            8'b01000010,
            8'b01111100,
            8'b01000000,
            8'b01000000,
            8'b01000000,
            8'b01000000
        };

        char[7'h52] = '{
            8'b01111100,
            8'b01000010,
            8'b01000010,
            8'b01111100,
            8'b01001000,
            8'b01000100,
            8'b01000010,
            8'b01000010
        };

        char[7'h53] = '{
            8'b00111100,
            8'b01000010,
            8'b01000000,
            8'b00111100,
            8'b00000010,
            8'b00000010,
            8'b01000010,
            8'b00111100
        };

        char[7'h54] = '{
            8'b01111110,
            8'b00011000,
            8'b00011000,
            8'b00011000,
            8'b00011000,
            8'b00011000,
            8'b00011000,
            8'b00011000
        };

        char[7'h56] = '{
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b00100100,
            8'b00011000,
            8'b00001000
        };

        char[7'h59] = '{
            8'b01000010,
            8'b01000010,
            8'b01000010,
            8'b00111100,
            8'b00011000,
            8'b00011000,
            8'b00011000,
            8'b00011000
        };
    end

    assign data = char[ascii_addr][char_row];

endmodule
